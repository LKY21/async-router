`timescale 1ns / 1ps
`include "macros.v"
`include "router.v"

module tree (CA4, CB4, CC5, CD5, CE6, CF6, CG7, CH7, C4A, C4B, C5C, C5D, C6E, C6F, C7G, C7H);
  
  `USES_CHANNEL
  parameter WIDTH = 11;
  
  `INPORT(CA4,WIDTH) 
  `INPORT(CB4,WIDTH) 
  `INPORT(CC5,WIDTH) 
  `INPORT(CD5,WIDTH) 
  `INPORT(CE6,WIDTH) 
  `INPORT(CF6,WIDTH) 
  `INPORT(CG7,WIDTH) 
  `INPORT(CH7,WIDTH) 

  `OUTPORT(C4A,WIDTH)
  `OUTPORT(C4B,WIDTH)  
  `OUTPORT(C5C,WIDTH)
  `OUTPORT(C5D,WIDTH)
  `OUTPORT(C6E,WIDTH)
  `OUTPORT(C6F,WIDTH)  
  `OUTPORT(C7G,WIDTH)
  `OUTPORT(C7H,WIDTH)  

  `CHANNEL(C10,WIDTH) 
  `CHANNEL(C01,WIDTH)
  `CHANNEL(C12,WIDTH) 
  `CHANNEL(C21,WIDTH)
  `CHANNEL(C24,WIDTH)
  `CHANNEL(C42,WIDTH)
  `CHANNEL(C25,WIDTH)
  `CHANNEL(C52,WIDTH)
  `CHANNEL(C4A,WIDTH)
  `CHANNEL(CA4,WIDTH)  
  `CHANNEL(C4B,WIDTH)
  `CHANNEL(CB4,WIDTH)
  `CHANNEL(C5C,WIDTH)
  `CHANNEL(CC5,WIDTH)
  `CHANNEL(C5D,WIDTH)
  `CHANNEL(CD5,WIDTH) 
  `CHANNEL(C13,WIDTH)
  `CHANNEL(C31,WIDTH)
  `CHANNEL(C36,WIDTH)
  `CHANNEL(C63,WIDTH)
  `CHANNEL(C37,WIDTH)
  `CHANNEL(C73,WIDTH)
  `CHANNEL(C6E,WIDTH) 
  `CHANNEL(CE6,WIDTH)
  `CHANNEL(C6F,WIDTH)
  `CHANNEL(CF6,WIDTH)
  `CHANNEL(C7G,WIDTH)
  `CHANNEL(CG7,WIDTH)
  `CHANNEL(C7H,WIDTH)  
  `CHANNEL(CH7,WIDTH)
    

  
//module router (C1, C2, P, C1out, C2out, Pout) ///oldd
 //module router (P, Pout, C1, C1out, C2, C2out)
 
  router R1(C01, C10, C21, C12, C31, C13);
  router R2(C12, C21, C42, C24, C52, C25);
  router R3(C13, C31, C63, C36, C73, C37);
  router R4(C24, C42, CA4, C4A, CB4, C4B);
  router R5(C25, C52, CC5, C5C, CD5, C5D);
  router R6(C36, C63, CE6, C6E, CF6, C6F);
  router R7(C37, C73, CG7, C7G, CH7, C7H);
endmodule
  
	
	
	
	
	
	
		

		
	

